* Generic MOS characterisation netlist

.param temp=27.000000
.temp 27.000000

* .lib "sky130_fd_pr/models/sky130.lib.spice" tt
.include "sky130_fd_pr/models/corners/tt.spice"

* circuit parameters
.param ids=1.200000
.param vds=1.800000
.param vdd=1.800000
.param vbs=1.200000
.param l=8.000000
.param vctl=-10

* the device under test
XM vd vg 0 vb sky130_fd_pr__pfet_01v8_mvt w=1 l=l m=1

* sources
Bgs 0 vg V=min(i(Vds)*1e9,vdd)
* BId 0 vd_ I=10**v(vctl)
Id vd_ 0 ids
Vds 0 vd_ DC={vds} AC=0
Vbs 0 vb {vbs}
Vctl vctl 0 {vctl}
Vdmeas vd_ vd
Hccvs out 0 Vdmeas 1

* specify op paramters to save
.save all @M.XM.msky130_fd_pr__pfet_01v8_mvt[id] @M.XM.msky130_fd_pr__pfet_01v8_mvt[vth] @M.XM.msky130_fd_pr__pfet_01v8_mvt[vgs] @M.XM.msky130_fd_pr__pfet_01v8_mvt[vds] @M.XM.msky130_fd_pr__pfet_01v8_mvt[vbs] @M.XM.msky130_fd_pr__pfet_01v8_mvt[gm] @M.XM.msky130_fd_pr__pfet_01v8_mvt[gds] @M.XM.msky130_fd_pr__pfet_01v8_mvt[gmbs] @M.XM.msky130_fd_pr__pfet_01v8_mvt[vdsat] @M.XM.msky130_fd_pr__pfet_01v8_mvt[cgg] @M.XM.msky130_fd_pr__pfet_01v8_mvt[cgs] @M.XM.msky130_fd_pr__pfet_01v8_mvt[cgd] @M.XM.msky130_fd_pr__pfet_01v8_mvt[cgb] @M.XM.msky130_fd_pr__pfet_01v8_mvt[cbs] @M.XM.msky130_fd_pr__pfet_01v8_mvt[cdd] 

* specify the simulations
.op
.noise v(out) Vds dec 10 1 1000Meg

* run the simulation and save the outputs
.control
  run
  setplot op1
  write spiceinterface_temp_op1.raw
  setplot noise1
  write spiceinterface_temp_noise1.raw
  quit
.endc

.end
